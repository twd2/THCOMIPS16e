library IEEE;
use IEEE.std_logic_1164.all;

package constants is
    constant ADDR_WIDTH: integer := 18;
    constant WORD_WIDTH: integer := 16;
end;